-- A DUT entity is used to wrap your design.
--  This example shows how you can do this for the
--  Full-adder.

library ieee;
use ieee.std_logic_1164.all;
entity DUT is
   port(input_vector: in std_logic_vector(2 downto 0);
       	output_vector: out std_logic_vector(0 downto 0));
end entity;

architecture DutWrap of DUT is
   component MUX  is
  port (A: in std_logic_vector(2 downto 0); O: out std_logic);
end component MUX;
begin

   -- input/output vector element ordering is critical,
   -- and must match the ordering in the trace file!
   add_instance: MUX 
			port map (
					-- order of inputs Cin B A
					A   => input_vector,                         -- order of outputs S Cout
					O => output_vector(0));

end DutWrap;

