-- A DUT entity is used to wrap your design.
--  This example shows how you can do this for the
--  Full-adder.

library ieee;
use ieee.std_logic_1164.all;
entity DUT is
   port(input_vector: in std_logic_vector(7 downto 0);
       	output_vector: out std_logic_vector(1 downto 0));
end entity;

architecture DutWrap of DUT is
   component Compare  is
  port (A: in std_logic_vector(7 downto 0);			
		  S:out std_logic_vector(1 downto 0));
end component Compare;
begin

   -- input/output vector element ordering is critical,
   -- and must match the ordering in the trace file!
   add_instance: Compare 
			port map (
					-- order of inputs Cin B A
					A   => input_vector,                         -- order of outputs S Cout
					S => output_vector);

end DutWrap;

